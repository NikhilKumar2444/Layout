*** SPICE deck for cell CMOS_inverter{lay} from library nikhil
*** Created on Mon May 19, 2025 22:46:01
*** Last revised on Thu May 22, 2025 23:05:20
*** Written on Thu May 22, 2025 23:05:33 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*** WARNING: no power connection for P-transistor wells in cell 'CMOS_inverter{lay}'
*** WARNING: no ground connection for N-transistor wells in cell 'CMOS_inverter{lay}'

*** TOP LEVEL CELL: CMOS_inverter{lay}
Mnmos@0 A_Not A nmos@0_diff-top gnd nmos_1 L=0.4U W=2.4U AS=1.44P AD=11.28P PS=6U PD=20.4U
Mpmos@0 A_Not A pmos@0_diff-top vdd pmos_1 L=0.4U W=2.4U AS=1.44P AD=11.28P PS=6U PD=20.4U

* Spice Code nodes in cell cell 'CMOS_inverter{lay}'
* CMOS Inverter Simulation in LTspice
* Power supply
Vdd Vdd 0 DC 5
* Input signal
Vin A 0 PULSE(0 5 10n 0.5n 0.5n 20n)
* Load capacitance
Cload A_Not 0 500f
* PMOS transistor (pull-up)
MpMOS A_Not A Vdd Vdd pmos_1 L=0.4u W=2.4u
* NMOS transistor (pull-down)
MnMOS A_Not A 0 0 nmos_1 L=0.4u W=2.4u
* Transistor models (renamed)
.model nmos_1 NMOS (LEVEL=1 VTO=0.7 KP=120u)
.model pmos_1 PMOS (LEVEL=1 VTO=-0.7 KP=50u)
* Transient simulation
.tran 0.1n 40n
.end
.END
