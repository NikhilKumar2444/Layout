*** SPICE deck for cell CMOS_nor{lay} from library nikhil
*** Created on Wed Jun 11, 2025 23:18:39
*** Last revised on Thu Jun 12, 2025 23:03:47
*** Written on Thu Jun 12, 2025 23:03:59 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: CMOS_nor{lay}
Mnmos@0 A_NOR_B A gnd gnd nMOS L=0.4U W=2.4U AS=5.52P AD=2.48P PS=13.2U PD=5.267U
Mnmos@2 gnd B A_NOR_B gnd nMOS L=0.4U W=2.4U AS=2.48P AD=5.52P PS=5.267U PD=13.2U
Mpmos@0 net@49 A vdd vdd pMOS L=0.4U W=2.4U AS=7.92P AD=1.62P PS=19U PD=6U
Mpmos@1 A_NOR_B B net@49 vdd pMOS L=0.4U W=2.4U AS=1.62P AD=2.48P PS=6U PD=5.267U

* Spice Code nodes in cell cell 'CMOS_nor{lay}'
* 2-input CMOS NAND Gate
* Inputs: A, B
* Output: A_NOR_B
* Power supply
Vdd vdd 0 DC 5
* Input signals
VinA A 0 PULSE(0 5 0ns 0.1ns 0.1ns 10ns 20ns)
VinB B 0 PULSE(0 5 0ns 0.1ns 0.1ns 20ns 40ns)
* Load at output
Cload A_NOR_B 0 500f
* PMOS pull-up network (parallel)
M1 A_NOR_B A vdd vdd pMOS L=0.4u W=2.4u
M2 A_NOR_B B vdd vdd pMOS L=0.4u W=2.4u
* NMOS pull-down network (series)
M3 net1 A 0 0 nMOS L=0.4u W=2.4u
M4 A_NOR_B B net1 0 nMOS L=0.4u W=2.4u
* Transistor models
.model nMOS NMOS (LEVEL=1 VTO=0.7 KP=120u)
.model pMOS PMOS (LEVEL=1 VTO=-0.7 KP=50u)
* Simulation command
.tran 0.1n 100n
.end
.END
