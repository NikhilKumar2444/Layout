*** SPICE deck for cell CMOS_nand{lay} from library nikhil
*** Created on Sun May 25, 2025 10:52:01
*** Last revised on Sun May 25, 2025 23:47:55
*** Written on Wed Jun 11, 2025 01:02:00 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: CMOS_nand{lay}
Mnmos@0 net@3 A gnd gnd nMOS L=0.4U W=2.4U AS=7.92P AD=1.2P PS=19U PD=3.4U
Mnmos@1 A_NAND_B B net@3 gnd nMOS L=0.4U W=2.4U AS=1.2P AD=2.48P PS=3.4U PD=5.267U
Mpmos@1 A_NAND_B A vdd vdd pMOS L=0.4U W=2.4U AS=5.52P AD=2.48P PS=13.2U PD=5.267U
Mpmos@3 vdd B A_NAND_B vdd pMOS L=0.4U W=2.4U AS=2.48P AD=5.52P PS=5.267U PD=13.2U

* Spice Code nodes in cell cell 'CMOS_nand{lay}'
* 2-input CMOS NAND Gate
* Inputs: A, B
* Output: A_NAND_B
* Power supply
Vdd vdd 0 DC 5
* Input signals
VinA A 0 PULSE(0 5 0ns 0.1ns 0.1ns 10ns 20ns)
VinB B 0 PULSE(0 5 0ns 0.1ns 0.1ns 20ns 40ns)
* Load at output
Cload A_NAND_B 0 500f
* PMOS pull-up network (parallel)
M1 A_NAND_B A vdd vdd pMOS L=0.4u W=2.4u
M2 A_NAND_B B vdd vdd pMOS L=0.4u W=2.4u
* NMOS pull-down network (series)
M3 net1 A 0 0 nMOS L=0.4u W=2.4u
M4 A_NAND_B B net1 0 nMOS L=0.4u W=2.4u
* Transistor models
.model nMOS NMOS (LEVEL=1 VTO=0.7 KP=120u)
.model pMOS PMOS (LEVEL=1 VTO=-0.7 KP=50u)
* Simulation command
.tran 0.1n 100n
.end
.END
